/**
 * Nand gate: 
 * out = 0 if (a == 1 and b == 1)
 *       1 otherwise
 */

 
module Nand(
	input a,
	input b,
	output out
);

	// No need to implement this chip
	// This chip is implemented using verilog primitives
	nand(out,a,b);

endmodule
