/**
* 9 bit Shiftregister (shifts to right)
* if      (load == 1)  out[t+1] = in[t]
* else if (shift == 1) out[t+1] = out[t]>>1 | (inMSB<<8)
* (shift one position to right and insert inMSB as most significant bit)
*/

 
module BitShift9R(
	input clk,
	input [8:0] in,
	input inMSB,
	input load,
	input shift,
	output [8:0] out
);

	// Put your code here:
	reg [8:0] shift_reg;
	always @(posedge clk) begin
		if (load == 1) begin
			shift_reg <= in;
		end else if (shift == 1) begin
			shift_reg <= (shift_reg  >> 1) | (inMSB<<8);
		end
	end
	assign out = shift_reg;

endmodule
